library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

package lpc_vectors is
    type lpc_interface is record
        lframe: std_logic;
        lad: std_logic_vector(3 downto 0);
    end record;
    type LPC_TEST_DATA is array(natural range <>) of lpc_interface;
    constant lpc_io_read : LPC_TEST_DATA := (
        ('1', "0000"),
        ('1', "0000"),
        ('0', "0000"), -- START
        ('1', "0000"), -- CYCTYPE + DIR : IO Read
        ('1', "0000"), -- ADDR most significant nibble
        ('1', "0000"),
        ('1', "1000"),
        ('1', "0000"), -- ADDR lease significant nibble
        ('1', "1111"), -- TAR
        ('1', "0000"), -- TAR
        ('1', "0101"), -- SYNC Short Wait
        ('1', "0000"), -- SYNC Ready
        ('1', "1010"), -- DATA
        ('1', "0101"), -- DATA
        ('1', "1111"), -- TAR
        ('1', "0000") -- TAR
    );
    constant lpc_io_write : LPC_TEST_DATA := (
        ('1', "0000"),
        ('1', "0000"),
        ('0', "0000"), -- START
        ('1', "0010"), -- CYCTYPE + DIR : IO Write
        ('1', "0000"), -- ADDR most significant nibble
        ('1', "0000"),
        ('1', "1000"),
        ('1', "0000"), -- ADDR lease significant nibble
        ('1', "1010"), -- DATA
        ('1', "0101"), -- DATA
        ('1', "1111"), -- TAR
        ('1', "0000"), -- TAR
        ('1', "0000"), -- SYNC
        ('1', "1111"), -- TAR
        ('1', "0000") -- TAR
    );
    constant lpc_mem_read : LPC_TEST_DATA := (
        ('1', "0000"),
        ('1', "0000"),
        ('0', "0000"), -- START
        ('1', "0100"), -- CYCTYPE + DIR : Memory Read
        ('1', "0000"), -- ADDR most significant nibble
        ('1', "0001"),
        ('1', "0010"),
        ('1', "0011"),
        ('1', "0100"),
        ('1', "0101"),
        ('1', "0110"),
        ('1', "0111"), -- ADDR lease significant nibble
        ('1', "1111"), -- TAR
        ('1', "0000"), -- TAR
        ('1', "0110"), -- SYNC Long
        ('1', "0110"), -- SYNC Long
        ('1', "0110"), -- SYNC Long
        ('1', "0110"), -- SYNC Long
        ('1', "0000"), -- SYNC Ready
        ('1', "1010"), -- DATA
        ('1', "0101"), -- DATA
        ('1', "1111"), -- TAR
        ('1', "0000") -- TAR
    );
    
    constant lpc_mem_write : LPC_TEST_DATA := (
        ('1', "0000"),
        ('1', "0000"),
        ('0', "1110"), -- START
        ('0', "0000"), -- START
        ('1', "0110"), -- CYCTYPE + DIR : Memory Write
        ('1', "0000"), -- ADDR most significant nibble
        ('1', "0001"),
        ('1', "0010"),
        ('1', "0011"),
        ('1', "0100"),
        ('1', "0101"),
        ('1', "0110"),
        ('1', "0111"), -- ADDR lease significant nibble
        ('1', "1010"), -- DATA
        ('1', "0101"), -- DATA
        ('1', "1111"), -- TAR
        ('1', "0000"), -- TAR
        ('1', "0000"), -- SYNC Ready
        ('1', "1111"), -- TAR
        ('1', "0000") -- TAR
    );
    
    constant lpc_dma_r8 : LPC_TEST_DATA := (
        ('1', "0000"),
        ('1', "0000"),
        ('0', "0000"), -- START
        ('1', "1000"), -- CYCTYPE + DIR : DMA Read
        ('1', "0011"), -- CHANNEL
        ('1', "0000"), -- SIZE : 8 bit
        ('1', "1010"), -- DATA
        ('1', "0101"), -- DATA
        ('1', "1111"), -- TAR
        ('1', "0000"), -- TAR
        ('1', "1001"), -- SYNC Ready
        ('1', "1111"), -- TAR
        ('1', "0000") -- TAR
    );
    
    constant lpc_dma_r16 : LPC_TEST_DATA := (
        ('1', "0000"),
        ('1', "0000"),
        ('0', "0000"), -- START
        ('1', "1000"), -- CYCTYPE + DIR : DMA Read
        ('1', "0010"), -- CHANNEL
        ('1', "0001"), -- SIZE : 16 bit
        ('1', "1010"), -- DATA
        ('1', "0101"), -- DATA
        ('1', "1111"), -- TAR
        ('1', "0000"), -- TAR
        ('1', "1001"), -- SYNC Ready
        ('1', "1111"), -- TAR
        ('1', "0000"), -- TAR
        ('1', "1010"), -- DATA
        ('1', "0101"), -- DATA
        ('1', "1111"), -- TAR
        ('1', "0000"), -- TAR
        ('1', "1001"), -- SYNC Ready
        ('1', "1111"), -- TAR
        ('1', "0000") -- TAR
    );

    constant lpc_dma_r32 : LPC_TEST_DATA := (
        ('1', "0000"),
        ('1', "0000"),
        ('0', "0000"), -- START
        ('1', "1000"), -- CYCTYPE + DIR : DMA Read
        ('1', "0111"), -- CHANNEL
        ('1', "0011"), -- SIZE : 32 bit
        ('1', "1010"), -- DATA
        ('1', "0101"), -- DATA
        ('1', "1111"), -- TAR
        ('1', "0000"), -- TAR
        ('1', "1001"), -- SYNC Ready
        ('1', "1111"), -- TAR
        ('1', "0000"), -- TAR
        ('1', "1010"), -- DATA
        ('1', "0101"), -- DATA
        ('1', "1111"), -- TAR
        ('1', "0000"), -- TAR
        ('1', "1001"), -- SYNC Ready
        ('1', "1111"), -- TAR
        ('1', "0000"), -- TAR
        ('1', "1010"), -- DATA
        ('1', "0101"), -- DATA
        ('1', "1111"), -- TAR
        ('1', "0000"), -- TAR
        ('1', "1001"), -- SYNC Ready
        ('1', "1111"), -- TAR
        ('1', "0000"), -- TAR
        ('1', "1010"), -- DATA
        ('1', "0101"), -- DATA
        ('1', "1111"), -- TAR
        ('1', "0000"), -- TAR
        ('1', "0000"), -- SYNC Ready
        ('1', "1111"), -- TAR
        ('1', "0000") -- TAR
    );
    
    constant lpc_dma_w8 : LPC_TEST_DATA := (
        ('1', "0000"),
        ('1', "0000"),
        ('0', "0000"), -- START
        ('1', "1010"), -- CYCTYPE + DIR : DMA Write
        ('1', "0011"), -- CHANNEL
        ('1', "0000"), -- SIZE : 8 bit
        ('1', "1111"), -- TAR
        ('1', "0000"), -- TAR
        ('1', "1001"), -- SYNC Ready
        ('1', "1010"), -- DATA
        ('1', "0101"), -- DATA
        ('1', "1111"), -- TAR
        ('1', "0000") -- TAR
    );
    
    constant lpc_dma_w16 : LPC_TEST_DATA := (
        ('1', "0000"),
        ('1', "0000"),
        ('0', "0000"), -- START
        ('1', "1010"), -- CYCTYPE + DIR : DMA Write
        ('1', "0011"), -- CHANNEL
        ('1', "0001"), -- SIZE : 16 bit
        ('1', "1111"), -- TAR
        ('1', "0000"), -- TAR
        ('1', "1001"), -- SYNC Ready
        ('1', "1010"), -- DATA
        ('1', "0101"), -- DATA
        ('1', "1001"), -- SYNC Ready
        ('1', "1010"), -- DATA
        ('1', "0101"), -- DATA
        ('1', "1111"), -- TAR
        ('1', "0000") -- TAR
    );

    constant lpc_dma_w32 : LPC_TEST_DATA := (
        ('1', "0000"),
        ('1', "0000"),
        ('0', "0000"), -- START
        ('1', "1010"), -- CYCTYPE + DIR : DMA Write
        ('1', "0011"), -- CHANNEL
        ('1', "0011"), -- SIZE : 32 bit
        ('1', "1111"), -- TAR
        ('1', "0000"), -- TAR
        ('1', "1001"), -- SYNC Ready
        ('1', "1010"), -- DATA
        ('1', "0101"), -- DATA
        ('1', "1001"), -- SYNC Ready
        ('1', "1010"), -- DATA
        ('1', "0101"), -- DATA
        ('1', "1001"), -- SYNC Ready
        ('1', "1010"), -- DATA
        ('1', "0101"), -- DATA
        ('1', "1001"), -- SYNC Ready
        ('1', "1010"), -- DATA
        ('1', "0101"), -- DATA
        ('1', "1111"), -- TAR
        ('1', "0000") -- TAR
    );
    
    constant lpc_bm_io_r8 : LPC_TEST_DATA := (
        ('1', "0000"),
        ('1', "0000"),
        ('0', "0010"), -- START
        ('1', "1111"), -- TAR
        ('1', "0000"), -- TAR
        ('1', "0000"), -- CYCTYPE + DIR : IO Read
        ('1', "0000"), -- ADDR most significant nibble
        ('1', "0000"),
        ('1', "1000"),
        ('1', "0000"), -- ADDR lease significant nibble
        ('1', "0000"), -- SIZE : 8 bits
        ('1', "1111"), -- TAR
        ('1', "0000"), -- TAR
        ('1', "0101"), -- SYNC Short Wait
        ('1', "0000"), -- SYNC Ready
        ('1', "1010"), -- DATA
        ('1', "0101"), -- DATA
        ('1', "1111"), -- TAR
        ('1', "0000") -- TAR
    );
    
    constant lpc_bm_io_r16 : LPC_TEST_DATA := (
        ('1', "0000"),
        ('1', "0000"),
        ('0', "0011"), -- START
        ('1', "1111"), -- TAR
        ('1', "0000"), -- TAR
        ('1', "0000"), -- CYCTYPE + DIR : IO Read
        ('1', "0000"), -- ADDR most significant nibble
        ('1', "0000"),
        ('1', "1000"),
        ('1', "0000"), -- ADDR lease significant nibble
        ('1', "0001"), -- SIZE : 16 bits
        ('1', "1111"), -- TAR
        ('1', "0000"), -- TAR
        ('1', "0101"), -- SYNC Short Wait
        ('1', "0000"), -- SYNC Ready
        ('1', "1010"), -- DATA
        ('1', "0101"), -- DATA
        ('1', "1010"), -- DATA
        ('1', "0101"), -- DATA
        ('1', "1111"), -- TAR
        ('1', "0000") -- TAR
    );
    constant lpc_bm_io_r32 : LPC_TEST_DATA := (
        ('1', "0000"),
        ('1', "0000"),
        ('0', "0010"), -- START
        ('1', "1111"), -- TAR
        ('1', "0000"), -- TAR
        ('1', "0000"), -- CYCTYPE + DIR : IO Read
        ('1', "0000"), -- ADDR most significant nibble
        ('1', "0000"),
        ('1', "1000"),
        ('1', "0000"), -- ADDR lease significant nibble
        ('1', "0011"), -- SIZE : 32 bits
        ('1', "1111"), -- TAR
        ('1', "0000"), -- TAR
        ('1', "0101"), -- SYNC Short Wait
        ('1', "0000"), -- SYNC Ready
        ('1', "1010"), -- DATA
        ('1', "1010"), -- DATA
        ('1', "0101"), -- DATA
        ('1', "1010"), -- DATA
        ('1', "0101"), -- DATA
        ('1', "1010"), -- DATA
        ('1', "0101"), -- DATA
        ('1', "0101"), -- DATA
        ('1', "1111"), -- TAR
        ('1', "0000") -- TAR
    );
    
    constant lpc_bm_io_w8 : LPC_TEST_DATA := (
        ('1', "0000"),
        ('1', "0000"),
        ('0', "0010"), -- START
        ('1', "1111"), -- TAR
        ('1', "0000"), -- TAR
        ('1', "0010"), -- CYCTYPE + DIR : IO Write
        ('1', "0000"), -- ADDR most significant nibble
        ('1', "0000"),
        ('1', "1000"),
        ('1', "0000"), -- ADDR lease significant nibble
        ('1', "0000"), -- SIZE : 8 bits
        ('1', "1010"), -- DATA
        ('1', "0101"), -- DATA
        ('1', "1111"), -- TAR
        ('1', "0000"), -- TAR
        ('1', "0101"), -- SYNC Short Wait
        ('1', "0000"), -- SYNC Ready
        ('1', "1111"), -- TAR
        ('1', "0000") -- TAR
    );
    
    constant lpc_bm_io_w16 : LPC_TEST_DATA := (
        ('1', "0000"),
        ('1', "0000"),
        ('0', "0011"), -- START
        ('1', "1111"), -- TAR
        ('1', "0000"), -- TAR
        ('1', "0010"), -- CYCTYPE + DIR : IO Write
        ('1', "0000"), -- ADDR most significant nibble
        ('1', "0000"),
        ('1', "1000"),
        ('1', "0000"), -- ADDR lease significant nibble
        ('1', "0001"), -- SIZE : 16 bits
        ('1', "1010"), -- DATA
        ('1', "0101"), -- DATA
        ('1', "1010"), -- DATA
        ('1', "0101"), -- DATA
        ('1', "1111"), -- TAR
        ('1', "0000"), -- TAR
        ('1', "0101"), -- SYNC Short Wait
        ('1', "0000"), -- SYNC Ready
        ('1', "1111"), -- TAR
        ('1', "0000") -- TAR
    );
    constant lpc_bm_io_w32 : LPC_TEST_DATA := (
        ('1', "0000"),
        ('1', "0000"),
        ('0', "0010"), -- START
        ('1', "1111"), -- TAR
        ('1', "0000"), -- TAR
        ('1', "0010"), -- CYCTYPE + DIR : IO Write
        ('1', "0000"), -- ADDR most significant nibble
        ('1', "0000"),
        ('1', "1000"),
        ('1', "0000"), -- ADDR lease significant nibble
        ('1', "0011"), -- SIZE : 32 bits
        ('1', "1010"), -- DATA
        ('1', "1010"), -- DATA
        ('1', "0101"), -- DATA
        ('1', "1010"), -- DATA
        ('1', "0101"), -- DATA
        ('1', "1010"), -- DATA
        ('1', "0101"), -- DATA
        ('1', "0101"), -- DATA
        ('1', "1111"), -- TAR
        ('1', "0000"), -- TAR
        ('1', "0101"), -- SYNC Short Wait
        ('1', "0000"), -- SYNC Ready
        ('1', "1111"), -- TAR
        ('1', "0000") -- TAR
    );
    
    constant lpc_bm_mem_r8 : LPC_TEST_DATA := (
        ('1', "0000"),
        ('1', "0000"),
        ('0', "0010"), -- START
        ('1', "1111"), -- TAR
        ('1', "0000"), -- TAR
        ('1', "0100"), -- CYCTYPE + DIR : Mem Read
        ('1', "0000"), -- ADDR most significant nibble
        ('1', "0000"),
        ('1', "1000"),
        ('1', "0000"),
        ('1', "0000"),
        ('1', "0000"),
        ('1', "1000"),
        ('1', "0000"), -- ADDR lease significant nibble
        ('1', "0000"), -- SIZE : 8 bits
        ('1', "1111"), -- TAR
        ('1', "0000"), -- TAR
        ('1', "0101"), -- SYNC Short Wait
        ('1', "0000"), -- SYNC Ready
        ('1', "1010"), -- DATA
        ('1', "0101"), -- DATA
        ('1', "1111"), -- TAR
        ('1', "0000") -- TAR
    );
    
    constant lpc_bm_mem_r16 : LPC_TEST_DATA := (
        ('1', "0000"),
        ('1', "0000"),
        ('0', "0011"), -- START
        ('1', "1111"), -- TAR
        ('1', "0000"), -- TAR
        ('1', "0100"), -- CYCTYPE + DIR : Mem Read
        ('1', "0000"), -- ADDR most significant nibble
        ('1', "0000"),
        ('1', "1000"),
        ('1', "0000"),
        ('1', "0000"),
        ('1', "0000"),
        ('1', "1000"),
        ('1', "0000"), -- ADDR lease significant nibble
        ('1', "0001"), -- SIZE : 16 bits
        ('1', "1111"), -- TAR
        ('1', "0000"), -- TAR
        ('1', "0101"), -- SYNC Short Wait
        ('1', "0000"), -- SYNC Ready
        ('1', "1010"), -- DATA
        ('1', "0101"), -- DATA
        ('1', "1010"), -- DATA
        ('1', "0101"), -- DATA
        ('1', "1111"), -- TAR
        ('1', "0000") -- TAR
    );
    constant lpc_bm_mem_r32 : LPC_TEST_DATA := (
        ('1', "0000"),
        ('1', "0000"),
        ('0', "0010"), -- START
        ('1', "1111"), -- TAR
        ('1', "0000"), -- TAR
        ('1', "0100"), -- CYCTYPE + DIR : Mem Read
        ('1', "0000"), -- ADDR most significant nibble
        ('1', "0000"),
        ('1', "1000"),
        ('1', "0000"), 
        ('1', "0000"), 
        ('1', "0000"),
        ('1', "1000"),
        ('1', "0000"), -- ADDR lease significant nibble
        ('1', "0011"), -- SIZE : 32 bits
        ('1', "1111"), -- TAR
        ('1', "0000"), -- TAR
        ('1', "0101"), -- SYNC Short Wait
        ('1', "0000"), -- SYNC Ready
        ('1', "1010"), -- DATA
        ('1', "1010"), -- DATA
        ('1', "0101"), -- DATA
        ('1', "1010"), -- DATA
        ('1', "0101"), -- DATA
        ('1', "1010"), -- DATA
        ('1', "0101"), -- DATA
        ('1', "0101"), -- DATA
        ('1', "1111"), -- TAR
        ('1', "0000") -- TAR
    );
    
    constant lpc_bm_mem_w8 : LPC_TEST_DATA := (
        ('1', "0000"),
        ('1', "0000"),
        ('0', "0010"), -- START
        ('1', "1111"), -- TAR
        ('1', "0000"), -- TAR
        ('1', "0110"), -- CYCTYPE + DIR : Mem Write
        ('1', "0000"), -- ADDR most significant nibble
        ('1', "0000"),
        ('1', "1000"),
        ('1', "0000"), 
        ('1', "0000"), 
        ('1', "0000"),
        ('1', "1000"),
        ('1', "0000"), -- ADDR lease significant nibble
        ('1', "0000"), -- SIZE : 8 bits
        ('1', "1010"), -- DATA
        ('1', "0101"), -- DATA
        ('1', "1111"), -- TAR
        ('1', "0000"), -- TAR
        ('1', "0101"), -- SYNC Short Wait
        ('1', "0000"), -- SYNC Ready
        ('1', "1111"), -- TAR
        ('1', "0000") -- TAR
    );
    
    constant lpc_bm_mem_w16 : LPC_TEST_DATA := (
        ('1', "0000"),
        ('1', "0000"),
        ('0', "0011"), -- START
        ('1', "1111"), -- TAR
        ('1', "0000"), -- TAR
        ('1', "0110"), -- CYCTYPE + DIR : Mem Write
        ('1', "0000"), -- ADDR most significant nibble
        ('1', "0000"),
        ('1', "1000"),
        ('1', "0000"), 
        ('1', "0000"), 
        ('1', "0000"),
        ('1', "1000"),
        ('1', "0000"), -- ADDR lease significant nibble
        ('1', "0001"), -- SIZE : 16 bits
        ('1', "1010"), -- DATA
        ('1', "0101"), -- DATA
        ('1', "1010"), -- DATA
        ('1', "0101"), -- DATA
        ('1', "1111"), -- TAR
        ('1', "0000"), -- TAR
        ('1', "0101"), -- SYNC Short Wait
        ('1', "0000"), -- SYNC Ready
        ('1', "1111"), -- TAR
        ('1', "0000") -- TAR
    );
    constant lpc_bm_mem_w32 : LPC_TEST_DATA := (
        ('1', "0000"),
        ('1', "0000"),
        ('0', "0010"), -- START
        ('1', "1111"), -- TAR
        ('1', "0000"), -- TAR
        ('1', "0110"), -- CYCTYPE + DIR : IO Write
        ('1', "0000"), -- ADDR most significant nibble
        ('1', "0000"),
        ('1', "1000"),
        ('1', "0000"), 
        ('1', "0000"), 
        ('1', "0000"),
        ('1', "1000"),
        ('1', "0000"), -- ADDR lease significant nibble
        ('1', "0011"), -- SIZE : 32 bits
        ('1', "1010"), -- DATA
        ('1', "1010"), -- DATA
        ('1', "0101"), -- DATA
        ('1', "1010"), -- DATA
        ('1', "0101"), -- DATA
        ('1', "1010"), -- DATA
        ('1', "0101"), -- DATA
        ('1', "0101"), -- DATA
        ('1', "1111"), -- TAR
        ('1', "0000"), -- TAR
        ('1', "0101"), -- SYNC Short Wait
        ('1', "0000"), -- SYNC Ready
        ('1', "1111"), -- TAR
        ('1', "0000") -- TAR
    );
    constant fwh_r8 : LPC_TEST_DATA := (
        ('1', "0000"),
        ('1', "0000"),
        ('0', "1101"), -- START
        ('1', "0000"), -- IDSEL
        ('1', "0001"), -- ADDR most significant nibble
        ('1', "0010"),
        ('1', "0011"),
        ('1', "0100"),
        ('1', "0101"),
        ('1', "0110"),
        ('1', "0111"), -- ADDR lease significant nibble
        ('1', "0000"), -- MSIZE: 1 byte
        ('1', "1111"), -- TAR
        ('1', "1111"), -- TAR
        ('1', "1111"), -- SYNC Long
        ('1', "1111"), -- SYNC Long
        ('1', "1111"), -- SYNC Long
        ('1', "1111"), -- SYNC Long
        ('0', "1111"), -- SYNC Ready
        ('0', "1111"), -- DATA
        ('0', "1111"), -- DATA
        ('0', "1111"), -- TAR
        ('1', "1111") -- TAR
    );
    constant ec_command : LPC_TEST_DATA := (
        ('1', "0000"),
        ('1', "0000"),
        ('0', "0000"), -- START
        ('1', "0010"), -- CYCTYPE + DIR : IO Write
        ('1', "0000"), -- ADDR most significant nibble
        ('1', "1001"),
        ('1', "0001"),
        ('1', "0000"), -- ADDR lease significant nibble
        ('1', "0000"), -- DATA
        ('1', "0000"), -- DATA
        ('1', "1111"), -- TAR
        ('1', "1111"), -- TAR
        ('1', "0000"), -- SYNC
        ('1', "1111"), -- TAR
        ('1', "1111"), -- TAR
        ('1', "0000"),
        ('1', "0000"),
        ('0', "0000"), -- START
        ('1', "0010"), -- CYCTYPE + DIR : IO Write
        ('1', "0000"), -- ADDR most significant nibble
        ('1', "1001"),
        ('1', "0001"),
        ('1', "0001"), -- ADDR lease significant nibble
        ('1', "0010"), -- DATA
        ('1', "1100"), -- DATA
        ('1', "1111"), -- TAR
        ('1', "1111"), -- TAR
        ('1', "0000"), -- SYNC
        ('1', "1111"), -- TAR
        ('1', "1111") -- TAR
    );
    constant ec_wait : LPC_TEST_DATA := (
        ('1', "1111"),
        ('1', "1111"),
        ('0', "0000"), -- START
        ('1', "0010"), -- CYCTYPE + DIR : IO Write
        ('1', "0000"), -- ADDR most significant nibble
        ('1', "1001"),
        ('1', "0001"),
        ('1', "0000"), -- ADDR lease significant nibble
        ('1', "0000"), -- DATA
        ('1', "0000"), -- DATA
        ('1', "1111"), -- TAR
        ('1', "1111"), -- TAR
        ('1', "0000"), -- SYNC
        ('1', "1111"), -- TAR
        ('1', "1111"), -- TAR
        ('1', "1111"),
        ('1', "1111"),
        ('0', "0000"), -- START
        ('1', "0000"), -- CYCTYPE + DIR : IO Read
        ('1', "0000"), -- ADDR most significant nibble
        ('1', "1001"),
        ('1', "0001"),
        ('1', "0001"), -- ADDR lease significant nibble
        ('1', "1111"), -- TAR
        ('1', "1111"), -- TAR
        ('1', "0101"), -- SYNC Short Wait
        ('1', "0000"), -- SYNC Ready
        ('1', "0010"), -- DATA
        ('1', "1100"), -- DATA
        ('1', "1111"), -- TAR
        ('1', "1111") -- TAR
    );
    constant ec_done : LPC_TEST_DATA := (
        ('1', "0000"),
        ('1', "0000"),
        ('0', "0000"), -- START
        ('1', "0010"), -- CYCTYPE + DIR : IO Write
        ('1', "0000"), -- ADDR most significant nibble
        ('1', "1001"),
        ('1', "0001"),
        ('1', "0000"), -- ADDR lease significant nibble
        ('1', "0000"), -- DATA
        ('1', "0000"), -- DATA
        ('1', "1111"), -- TAR
        ('1', "1111"), -- TAR
        ('1', "0000"), -- SYNC
        ('1', "1111"), -- TAR
        ('1', "1111"), -- TAR
        ('1', "0000"),
        ('1', "0000"),
        ('0', "0000"), -- START
        ('1', "0000"), -- CYCTYPE + DIR : IO Read
        ('1', "0000"), -- ADDR most significant nibble
        ('1', "1001"),
        ('1', "0001"),
        ('1', "0001"), -- ADDR lease significant nibble
        ('1', "1111"), -- TAR
        ('1', "1111"), -- TAR
        ('1', "0101"), -- SYNC Short Wait
        ('1', "0000"), -- SYNC Ready
        ('1', "0000"), -- DATA
        ('1', "0000"), -- DATA
        ('1', "1111"), -- TAR
        ('1', "1111") -- TAR
    );
    constant lpc_io_84_write : LPC_TEST_DATA := (
        ('1', "0000"),
        ('1', "0000"),
        ('0', "0000"), -- START
        ('1', "0010"), -- CYCTYPE + DIR : IO Write
        ('1', "0000"), -- ADDR most significant nibble
        ('1', "0000"),
        ('1', "1000"),
        ('1', "0100"), -- ADDR lease significant nibble
        ('1', "0001"), -- DATA
        ('1', "0100"), -- DATA
        ('1', "1111"), -- TAR
        ('1', "1111"), -- TAR
        ('1', "1111"), -- SYNC
        ('1', "1111"), -- SYNC
        ('1', "1111"), -- SYNC
        ('1', "1111"), -- SYNC
        ('0', "1111"), -- TAR
        ('0', "1111"), -- TAR
        ('0', "1111"), -- TAR
        ('0', "1111"), -- TAR
        ('1', "1111"), -- IDLE
        ('1', "1111") -- IDLE
    );
    constant e6400_test : LPC_TEST_DATA := ( 
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('0', "0000"),
        ('1', "0010"),
        ('1', "0000"),
        ('1', "0000"),
        ('1', "0010"),
        ('1', "1110"),
        ('1', "0101"),
        ('1', "0101"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "0110"),
        ('1', "0110"),
        ('1', "0110"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('0', "0000"),
        ('1', "0010"),
        ('1', "0000"),
        ('1', "0000"),
        ('1', "0010"),
        ('1', "1110"),
        ('1', "0101"),
        ('1', "0101"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "0110"),
        ('1', "0110"),
        ('1', "0110"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('0', "0000"),
        ('1', "0010"),
        ('1', "0000"),
        ('1', "0000"),
        ('1', "0010"),
        ('1', "1110"),
        ('1', "0100"),
        ('1', "0010"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "0110"),
        ('1', "0110"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('0', "0000"),
        ('1', "0010"),
        ('1', "0000"),
        ('1', "0000"),
        ('1', "0010"),
        ('1', "1111"),
        ('1', "0100"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "0110"),
        ('1', "0110"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('0', "0000"),
        ('1', "0010"),
        ('1', "0000"),
        ('1', "0000"),
        ('1', "0010"),
        ('1', "1110"),
        ('1', "1010"),
        ('1', "1010"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "0110"),
        ('1', "0110"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('0', "0000"),
        ('1', "0010"),
        ('1', "0000"),
        ('1', "1001"),
        ('1', "0100"),
        ('1', "1110"),
        ('1', "0101"),
        ('1', "0101"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "0110"),
        ('1', "0110"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('0', "0000"),
        ('1', "0010"),
        ('1', "0000"),
        ('1', "1001"),
        ('1', "0100"),
        ('1', "1110"),
        ('1', "0101"),
        ('1', "0101"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "0110"),
        ('1', "0110"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('0', "0000"),
        ('1', "0010"),
        ('1', "0000"),
        ('1', "1001"),
        ('1', "0100"),
        ('1', "1110"),
        ('1', "0010"),
        ('1', "0010"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "0110"),
        ('1', "0110"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('0', "0000"),
        ('1', "0010"),
        ('1', "0000"),
        ('1', "1001"),
        ('1', "0100"),
        ('1', "1111"),
        ('1', "0000"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "0110"),
        ('1', "0110"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('0', "0000"),
        ('1', "0010"),
        ('1', "0000"),
        ('1', "1001"),
        ('1', "0100"),
        ('1', "1110"),
        ('1', "0011"),
        ('1', "0010"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "0110"),
        ('1', "0110"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('0', "0000"),
        ('1', "0010"),
        ('1', "0000"),
        ('1', "1001"),
        ('1', "0100"),
        ('1', "1111"),
        ('1', "0000"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "0110"),
        ('1', "0110"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('0', "0000"),
        ('1', "0010"),
        ('1', "0000"),
        ('1', "1001"),
        ('1', "0100"),
        ('1', "1110"),
        ('1', "0100"),
        ('1', "0010"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "0110"),
        ('1', "0110"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('0', "0000"),
        ('1', "0010"),
        ('1', "0000"),
        ('1', "1001"),
        ('1', "0100"),
        ('1', "1111"),
        ('1', "0100"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "0110"),
        ('1', "0110"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('0', "0000"),
        ('1', "0010"),
        ('1', "0000"),
        ('1', "1001"),
        ('1', "0100"),
        ('1', "1110"),
        ('1', "0101"),
        ('1', "0010"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "0110"),
        ('1', "0110"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('0', "0000"),
        ('1', "0010"),
        ('1', "0000"),
        ('1', "1001"),
        ('1', "0100"),
        ('1', "1111"),
        ('1', "0100"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "0110"),
        ('1', "0110"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('0', "0000"),
        ('1', "0010"),
        ('1', "0000"),
        ('1', "1001"),
        ('1', "0100"),
        ('1', "1110"),
        ('1', "0111"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "0110"),
        ('1', "0110"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('0', "0000"),
        ('1', "0010"),
        ('1', "0000"),
        ('1', "1001"),
        ('1', "0100"),
        ('1', "1111"),
        ('1', "0011"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "0110"),
        ('1', "0110"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('0', "0000"),
        ('1', "0010"),
        ('1', "0000"),
        ('1', "1001"),
        ('1', "0100"),
        ('1', "1110"),
        ('1', "0000"),
        ('1', "0011"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "0110"),
        ('1', "0110"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('0', "0000"),
        ('1', "0010"),
        ('1', "0000"),
        ('1', "1001"),
        ('1', "0100"),
        ('1', "1111"),
        ('1', "0001"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "0110"),
        ('1', "0110"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('0', "0000"),
        ('1', "0010"),
        ('1', "0000"),
        ('1', "1001"),
        ('1', "0100"),
        ('1', "1110"),
        ('1', "0000"),
        ('1', "0110"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "0110"),
        ('1', "0110"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('0', "0000"),
        ('1', "0010"),
        ('1', "0000"),
        ('1', "1001"),
        ('1', "0100"),
        ('1', "1111"),
        ('1', "0000"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "0110"),
        ('1', "0110"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('0', "0000"),
        ('1', "0010"),
        ('1', "0000"),
        ('1', "1001"),
        ('1', "0100"),
        ('1', "1110"),
        ('1', "0001"),
        ('1', "0110"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "0110"),
        ('1', "0110"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('0', "0000"),
        ('1', "0010"),
        ('1', "0000"),
        ('1', "1001"),
        ('1', "0100"),
        ('1', "1111"),
        ('1', "0000"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "0110"),
        ('1', "0110"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('0', "0000"),
        ('1', "0010"),
        ('1', "0000"),
        ('1', "1001"),
        ('1', "0100"),
        ('1', "1110"),
        ('1', "0000"),
        ('1', "0111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "0110"),
        ('1', "0110"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('0', "0000"),
        ('1', "0010"),
        ('1', "0000"),
        ('1', "1001"),
        ('1', "0100"),
        ('1', "1111"),
        ('1', "0000"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "0110"),
        ('1', "0110"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('0', "0000"),
        ('1', "0010"),
        ('1', "0000"),
        ('1', "1001"),
        ('1', "0100"),
        ('1', "1110"),
        ('1', "0010"),
        ('1', "0111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "0110"),
        ('1', "0110"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('0', "0000"),
        ('1', "0010"),
        ('1', "0000"),
        ('1', "1001"),
        ('1', "0100"),
        ('1', "1111"),
        ('1', "0000"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "0110"),
        ('1', "0110"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('0', "0000"),
        ('1', "0010"),
        ('1', "0000"),
        ('1', "1001"),
        ('1', "0100"),
        ('1', "1110"),
        ('1', "0100"),
        ('1', "0111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "0110"),
        ('1', "0110"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('0', "0000"),
        ('1', "0010"),
        ('1', "0000"),
        ('1', "1001"),
        ('1', "0100"),
        ('1', "1111"),
        ('1', "0100"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "0110"),
        ('1', "0110"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('0', "0000"),
        ('1', "0010"),
        ('1', "0000"),
        ('1', "1001"),
        ('1', "0100"),
        ('1', "1110"),
        ('1', "0000"),
        ('1', "0011"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "0110"),
        ('1', "0110"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('0', "0000"),
        ('1', "0010"),
        ('1', "0000"),
        ('1', "1001"),
        ('1', "0100"),
        ('1', "1111"),
        ('1', "0001"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "0110"),
        ('1', "0110"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('0', "0000"),
        ('1', "0010"),
        ('1', "0000"),
        ('1', "1001"),
        ('1', "0100"),
        ('1', "1110"),
        ('1', "0000"),
        ('1', "0011"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "0110"),
        ('1', "0110"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('0', "0000"),
        ('1', "0010"),
        ('1', "0000"),
        ('1', "1001"),
        ('1', "0100"),
        ('1', "1111"),
        ('1', "0000"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "0110"),
        ('1', "0110"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('0', "0000"),
        ('1', "0010"),
        ('1', "0000"),
        ('1', "1001"),
        ('1', "0100"),
        ('1', "1110"),
        ('1', "0111"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "0110"),
        ('1', "0110"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('0', "0000"),
        ('1', "0010"),
        ('1', "0000"),
        ('1', "1001"),
        ('1', "0100"),
        ('1', "1111"),
        ('1', "0100"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "0110"),
        ('1', "0110"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('0', "0000"),
        ('1', "0010"),
        ('1', "0000"),
        ('1', "1001"),
        ('1', "0100"),
        ('1', "1110"),
        ('1', "0000"),
        ('1', "0011"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "0110"),
        ('1', "0110"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('0', "0000"),
        ('1', "0010"),
        ('1', "0000"),
        ('1', "1001"),
        ('1', "0100"),
        ('1', "1111"),
        ('1', "0001"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "0110"),
        ('1', "0110"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('0', "0000"),
        ('1', "0010"),
        ('1', "0000"),
        ('1', "1001"),
        ('1', "0100"),
        ('1', "1110"),
        ('1', "0000"),
        ('1', "0110"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "0110"),
        ('1', "0110"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('0', "0000"),
        ('1', "0010"),
        ('1', "0000"),
        ('1', "1001"),
        ('1', "0100"),
        ('1', "1111"),
        ('1', "0000"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "0110"),
        ('1', "0110"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('0', "0000"),
        ('1', "0010"),
        ('1', "0000"),
        ('1', "1001"),
        ('1', "0100"),
        ('1', "1110"),
        ('1', "0001"),
        ('1', "0110"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "0110"),
        ('1', "0110"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('0', "0000"),
        ('1', "0010"),
        ('1', "0000"),
        ('1', "1001"),
        ('1', "0100"),
        ('1', "1111"),
        ('1', "0000"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "0110"),
        ('1', "0110"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('0', "0000"),
        ('1', "0010"),
        ('1', "0000"),
        ('1', "1001"),
        ('1', "0100"),
        ('1', "1110"),
        ('1', "0000"),
        ('1', "0111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "0110"),
        ('1', "0110"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('0', "0000"),
        ('1', "0010"),
        ('1', "0000"),
        ('1', "1001"),
        ('1', "0100"),
        ('1', "1111"),
        ('1', "0000"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "0110"),
        ('1', "0110"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('0', "0000"),
        ('1', "0010"),
        ('1', "0000"),
        ('1', "1001"),
        ('1', "0100"),
        ('1', "1110"),
        ('1', "0010"),
        ('1', "0111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "0110"),
        ('1', "0110"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('0', "0000"),
        ('1', "0010"),
        ('1', "0000"),
        ('1', "1001"),
        ('1', "0100"),
        ('1', "1111"),
        ('1', "0000"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "0110"),
        ('1', "0110"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('0', "0000"),
        ('1', "0010"),
        ('1', "0000"),
        ('1', "1001"),
        ('1', "0100"),
        ('1', "1110"),
        ('1', "0000"),
        ('1', "0011"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "0110"),
        ('1', "0110"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('0', "0000"),
        ('1', "0010"),
        ('1', "0000"),
        ('1', "1001"),
        ('1', "0100"),
        ('1', "1111"),
        ('1', "0001"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "0110"),
        ('1', "0110"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('0', "0000"),
        ('1', "0010"),
        ('1', "0000"),
        ('1', "1001"),
        ('1', "0100"),
        ('1', "1110"),
        ('1', "0000"),
        ('1', "0011"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "0110"),
        ('1', "0110"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('0', "0000"),
        ('1', "0010"),
        ('1', "0000"),
        ('1', "1001"),
        ('1', "0100"),
        ('1', "1111"),
        ('1', "0000"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "0110"),
        ('1', "0110"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('0', "0000"),
        ('1', "0010"),
        ('1', "0000"),
        ('1', "1001"),
        ('1', "0100"),
        ('1', "1110"),
        ('1', "0111"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "0110"),
        ('1', "0110"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('0', "0000"),
        ('1', "0010"),
        ('1', "0000"),
        ('1', "1001"),
        ('1', "0100"),
        ('1', "1111"),
        ('1', "0101"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "0110"),
        ('1', "0110"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('0', "0000"),
        ('1', "0010"),
        ('1', "0000"),
        ('1', "1001"),
        ('1', "0100"),
        ('1', "1110"),
        ('1', "0000"),
        ('1', "0011"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "0110"),
        ('1', "0110"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('0', "0000"),
        ('1', "0010"),
        ('1', "0000"),
        ('1', "1001"),
        ('1', "0100"),
        ('1', "1111"),
        ('1', "0001"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "0110"),
        ('1', "0110"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('0', "0000"),
        ('1', "0010"),
        ('1', "0000"),
        ('1', "1001"),
        ('1', "0100"),
        ('1', "1110"),
        ('1', "0000"),
        ('1', "0110"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "0110"),
        ('1', "0110"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('0', "0000"),
        ('1', "0010"),
        ('1', "0000"),
        ('1', "1001"),
        ('1', "0100"),
        ('1', "1111"),
        ('1', "0000"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "0110"),
        ('1', "0110"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('0', "0000"),
        ('1', "0010"),
        ('1', "0000"),
        ('1', "1001"),
        ('1', "0100"),
        ('1', "1110"),
        ('1', "0001"),
        ('1', "0110"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "0110"),
        ('1', "0110"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('0', "0000"),
        ('1', "0010"),
        ('1', "0000"),
        ('1', "1001"),
        ('1', "0100"),
        ('1', "1111"),
        ('1', "0000"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "0110"),
        ('1', "0110"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('0', "0000"),
        ('1', "0010"),
        ('1', "0000"),
        ('1', "1001"),
        ('1', "0100"),
        ('1', "1110"),
        ('1', "0000"),
        ('1', "0111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "0110"),
        ('1', "0110"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('0', "0000"),
        ('1', "0010"),
        ('1', "0000"),
        ('1', "1001"),
        ('1', "0100"),
        ('1', "1111"),
        ('1', "0000"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "0110"),
        ('1', "0110"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('0', "0000"),
        ('1', "0010"),
        ('1', "0000"),
        ('1', "1001"),
        ('1', "0100"),
        ('1', "1110"),
        ('1', "0010"),
        ('1', "0111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "0110"),
        ('1', "0110"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('0', "0000"),
        ('1', "0010"),
        ('1', "0000"),
        ('1', "1001"),
        ('1', "0100"),
        ('1', "1111"),
        ('1', "0000"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "0110"),
        ('1', "0110"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('0', "0000"),
        ('1', "0010"),
        ('1', "0000"),
        ('1', "1001"),
        ('1', "0100"),
        ('1', "1110"),
        ('1', "0100"),
        ('1', "0111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "0110"),
        ('1', "0110"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('0', "0000"),
        ('1', "0010"),
        ('1', "0000"),
        ('1', "1001"),
        ('1', "0100"),
        ('1', "1111"),
        ('1', "0100"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "0110"),
        ('1', "0110"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('0', "0000"),
        ('1', "0010"),
        ('1', "0000"),
        ('1', "1001"),
        ('1', "0100"),
        ('1', "1110"),
        ('1', "0000"),
        ('1', "0011"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "0110"),
        ('1', "0110"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('0', "0000"),
        ('1', "0010"),
        ('1', "0000"),
        ('1', "1001"),
        ('1', "0100"),
        ('1', "1111"),
        ('1', "0001"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "0110"),
        ('1', "0110"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('0', "0000"),
        ('1', "0010"),
        ('1', "0000"),
        ('1', "1001"),
        ('1', "0100"),
        ('1', "1110"),
        ('1', "0000"),
        ('1', "0011"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "0110"),
        ('1', "0110"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('0', "0000"),
        ('1', "0010"),
        ('1', "0000"),
        ('1', "1001"),
        ('1', "0100"),
        ('1', "1111"),
        ('1', "0000"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "0110"),
        ('1', "0110"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('0', "0000"),
        ('1', "0010"),
        ('1', "0000"),
        ('1', "1001"),
        ('1', "0100"),
        ('1', "1110"),
        ('1', "0111"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "0110"),
        ('1', "0110"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('0', "0000"),
        ('1', "0010"),
        ('1', "0000"),
        ('1', "1001"),
        ('1', "0100"),
        ('1', "1111"),
        ('1', "1100"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "0110"),
        ('1', "0110"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('0', "0000"),
        ('1', "0010"),
        ('1', "0000"),
        ('1', "1001"),
        ('1', "0100"),
        ('1', "1110"),
        ('1', "0000"),
        ('1', "0011"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "0110"),
        ('1', "0110"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('0', "0000"),
        ('1', "0010"),
        ('1', "0000"),
        ('1', "1001"),
        ('1', "0100"),
        ('1', "1111"),
        ('1', "0001"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "0110"),
        ('1', "0110"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('0', "0000"),
        ('1', "0010"),
        ('1', "0000"),
        ('1', "1001"),
        ('1', "0100"),
        ('1', "1110"),
        ('1', "0000"),
        ('1', "0110"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "0110"),
        ('1', "0110"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('0', "0000"),
        ('1', "0010"),
        ('1', "0000"),
        ('1', "1001"),
        ('1', "0100"),
        ('1', "1111"),
        ('1', "1001"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "0110"),
        ('1', "0110"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('0', "0000"),
        ('1', "0010"),
        ('1', "0000"),
        ('1', "1001"),
        ('1', "0100"),
        ('1', "1110"),
        ('1', "0001"),
        ('1', "0110"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "0110"),
        ('1', "0110"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('0', "0000"),
        ('1', "0010"),
        ('1', "0000"),
        ('1', "1001"),
        ('1', "0100"),
        ('1', "1111"),
        ('1', "1000"),
        ('1', "0010"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "0110"),
        ('1', "0110"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('0', "0000"),
        ('1', "0010"),
        ('1', "0000"),
        ('1', "1001"),
        ('1', "0100"),
        ('1', "1110"),
        ('1', "0000"),
        ('1', "0111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "0110"),
        ('1', "0110"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('0', "0000"),
        ('1', "0010"),
        ('1', "0000"),
        ('1', "1001"),
        ('1', "0100"),
        ('1', "1111"),
        ('1', "0000"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "0110"),
        ('1', "0110"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('0', "0000"),
        ('1', "0010"),
        ('1', "0000"),
        ('1', "1001"),
        ('1', "0100"),
        ('1', "1110"),
        ('1', "0010"),
        ('1', "0111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "0110"),
        ('1', "0110"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('0', "0000"),
        ('1', "0010"),
        ('1', "0000"),
        ('1', "1001"),
        ('1', "0100"),
        ('1', "1111"),
        ('1', "0000"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "0110"),
        ('1', "0110"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('0', "0000"),
        ('1', "0010"),
        ('1', "0000"),
        ('1', "1001"),
        ('1', "0100"),
        ('1', "1110"),
        ('1', "0100"),
        ('1', "0111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "0110"),
        ('1', "0110"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('0', "0000"),
        ('1', "0010"),
        ('1', "0000"),
        ('1', "1001"),
        ('1', "0100"),
        ('1', "1111"),
        ('1', "0001"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "0110"),
        ('1', "0110"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('0', "0000"),
        ('1', "0010"),
        ('1', "0000"),
        ('1', "1001"),
        ('1', "0100"),
        ('1', "1110"),
        ('1', "0000"),
        ('1', "0011"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "0110"),
        ('1', "0110"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('0', "0000"),
        ('1', "0010"),
        ('1', "0000"),
        ('1', "1001"),
        ('1', "0100"),
        ('1', "1111"),
        ('1', "0001"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "0110"),
        ('1', "0110"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('0', "0000"),
        ('1', "0010"),
        ('1', "0000"),
        ('1', "1001"),
        ('1', "0100"),
        ('1', "1110"),
        ('1', "1010"),
        ('1', "1010"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "0110"),
        ('1', "0110"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('0', "0000"),
        ('1', "0010"),
        ('1', "0000"),
        ('1', "1001"),
        ('1', "0001"),
        ('1', "0000"),
        ('1', "0000"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "0110"),
        ('1', "0110"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('0', "0000"),
        ('1', "0010"),
        ('1', "0000"),
        ('1', "1001"),
        ('1', "0001"),
        ('1', "0001"),
        ('1', "0001"),
        ('1', "1100"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "0110"),
        ('1', "0110"),
        ('1', "0110"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('0', "0000"),
        ('1', "0010"),
        ('1', "0000"),
        ('1', "1001"),
        ('1', "0001"),
        ('1', "0000"),
        ('1', "0000"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "0110"),
        ('1', "0110"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('0', "0000"),
        ('1', "0000"),
        ('1', "0000"),
        ('1', "1001"),
        ('1', "0001"),
        ('1', "0001"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "0110"),
        ('1', "0110"),
        ('1', "0110"),
        ('1', "0000"),
        ('1', "0001"),
        ('1', "1100"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "1111"),
        ('0', "0000"),
        ('1', "0010"),
        ('1', "0000"),
        ('1', "1001"),
        ('1', "0001"),
        ('1', "0000"),
        ('1', "0000"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111"),
        ('1', "0110"),
        ('1', "0110"),
        ('1', "0000"),
        ('1', "1111"),
        ('1', "1111")
    );
end package;
